magic
tech sky130A
timestamp 1694482379
<< nwell >>
rect -190 0 25 140
<< nmos >>
rect -60 -135 -45 -35
<< pmos >>
rect -60 20 -45 120
<< ndiff >>
rect -115 -50 -60 -35
rect -115 -120 -95 -50
rect -75 -120 -60 -50
rect -115 -135 -60 -120
rect -45 -50 5 -35
rect -45 -120 -30 -50
rect -10 -120 5 -50
rect -45 -135 5 -120
<< pdiff >>
rect -115 105 -60 120
rect -115 35 -95 105
rect -75 35 -60 105
rect -115 20 -60 35
rect -45 105 5 120
rect -45 35 -30 105
rect -10 35 5 105
rect -45 20 5 35
<< ndiffc >>
rect -95 -120 -75 -50
rect -30 -120 -10 -50
<< pdiffc >>
rect -95 35 -75 105
rect -30 35 -10 105
<< psubdiff >>
rect -170 -50 -115 -35
rect -170 -120 -155 -50
rect -135 -120 -115 -50
rect -170 -135 -115 -120
<< nsubdiff >>
rect -170 105 -115 120
rect -170 35 -155 105
rect -135 35 -115 105
rect -170 20 -115 35
<< psubdiffcont >>
rect -155 -120 -135 -50
<< nsubdiffcont >>
rect -155 35 -135 105
<< poly >>
rect -60 120 -45 135
rect -60 -35 -45 20
rect -60 -150 -45 -135
rect -85 -160 -45 -150
rect -85 -180 -75 -160
rect -55 -180 -45 -160
rect -85 -190 -45 -180
<< polycont >>
rect -75 -180 -55 -160
<< locali >>
rect -165 105 -65 115
rect -165 35 -155 105
rect -135 35 -95 105
rect -75 35 -65 105
rect -165 25 -65 35
rect -40 105 0 115
rect -40 35 -30 105
rect -10 35 0 105
rect -40 25 0 35
rect -20 -40 0 25
rect -165 -50 -65 -40
rect -165 -120 -155 -50
rect -135 -120 -95 -50
rect -75 -120 -65 -50
rect -165 -130 -65 -120
rect -40 -50 0 -40
rect -40 -120 -30 -50
rect -10 -120 0 -50
rect -40 -130 0 -120
rect -20 -150 0 -130
rect -185 -160 -45 -150
rect -185 -170 -75 -160
rect -85 -180 -75 -170
rect -55 -180 -45 -160
rect -20 -170 20 -150
rect -85 -190 -45 -180
<< viali >>
rect -155 35 -135 105
rect -95 35 -75 105
rect -155 -120 -135 -50
rect -95 -120 -75 -50
<< metal1 >>
rect -185 105 20 115
rect -185 35 -155 105
rect -135 35 -95 105
rect -75 35 20 105
rect -185 25 20 35
rect -185 -50 20 -40
rect -185 -120 -155 -50
rect -135 -120 -95 -50
rect -75 -120 20 -50
rect -185 -130 20 -120
<< labels >>
rlabel locali -185 -160 -185 -160 7 A
port 1 w
rlabel locali 20 -160 20 -160 3 Y
port 2 e
rlabel metal1 -185 70 -185 70 7 VP
port 3 w
rlabel metal1 -185 -85 -185 -85 7 VN
port 4 w
<< end >>

magic
tech sky130A
timestamp 1694482379
<< psubdiff >>
rect 0 0 55 85
<< ndiff >>
rect 55 0 170 85
<< poly >>
rect 105 -15 120 85
<< locali >>
rect 5 5 100 85
rect 125 5 165 85
<< ndiffc >>
rect 135 15 155 85
rect 20 15 40 85
rect 70 15 90 85
<< viali >>
rect 20 15 40 85
rect 70 15 90 85
<< metal1 >>
rect -15 5 185 85
<< nmos >>
rect 105 85 120 100
<< ndiff >>
rect 55 85 105 100
rect 120 85 170 100
<< psubdiff >>
rect 0 85 55 100
<< poly >>
rect 105 100 120 115
<< locali >>
rect 5 85 100 95
rect 125 85 165 95
<< metal1 >>
rect -15 85 185 95
<< end >>
